module simple_14 (
    input [4:0] a,
    input [4:0] b,
    output [3:0] sum
  );
    assign sum = a + b;
endmodule
