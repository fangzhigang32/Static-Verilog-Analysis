module medium_14 (
    input wire [3:0] a,
    input wire [3:0] b,
    output wire [7:0] sum
);
    assign sum = a + b;
endmodule
