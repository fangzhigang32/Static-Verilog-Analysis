module simple_30 (
    input wire a,
    input wire b,
    output reg c
  );
    assign c = a + b;
endmodule
