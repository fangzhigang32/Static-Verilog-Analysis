module simple_21(
    input a,
    input b,
    input cin,
    output sum
    );
    and (a,b,cin);
    assign sum = a;
endmodule