module medium_17(
    input a,
    output cout
);
    and (cout,a);
endmodule